interface shift_if(input clk);
    logic in;
    logic out;
endinterface : shift_if