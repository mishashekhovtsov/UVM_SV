interface shift_if(input clk, input rst_n);
    logic in;
    logic out;
    logic oe;
endinterface : shift_if