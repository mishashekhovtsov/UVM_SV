import uvm_pkg::*;
`include "uvm_macros.svh"

import shift_pkg::*;
import clk_gen_pkg::*;
import rst_gen_pkg::*;

`include "../uvm_classes/vseqr_cls.svh"
`include "../uvm_classes/base_vseq.svh"
`include "../uvm_classes/scb.svh"
`include "../uvm_classes/env.svh"
`include "../uvm_classes/base_test.svh"

