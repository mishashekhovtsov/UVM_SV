import uvm_pkg::*;
`include "uvm_macros.svh"

import shift_pkg::*;
import clk_gen_pkg::*;
import rst_gen_pkg::*;

`include "vseqr_cls.svh"
`include "scb.svh"
`include "env.svh"

`include "base_vseq.svh"
`include "SHIFT_VSEQ.svh"

`include "base_test.svh"
