interface shift_if(input clk, input rst_n);
    logic in;
    logic out;
endinterface : shift_if