package tb_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import shift_pkg::*;

    `include "../uvm_classes/shift_scb.svh"
    `include "../uvm_classes/env.svh"
    `include "../uvm_classes/base_test.svh"

endpackage : tb_pkg
